package frame_en_lib;
    `define hsv_v3                      1
endpackage
