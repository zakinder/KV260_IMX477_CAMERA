--01062019 [01-06-2019]
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.tbPackage.all;
use work.constants_package.all;
use work.vpf_records.all;
entity dut_configAxis is 
generic (
    aclk_freq                 : real    := 75.00e6;
    C_vfpConfig_DATA_WIDTH    : integer := 32;
    C_vfpconfig_ADDR_WIDTH    : integer := 8);
port (
    vfpconfig_aclk            : out std_logic;
    vfpconfig_aresetn         : out std_logic;
    vfpconfig_awaddr          : out std_logic_vector(C_vfpconfig_ADDR_WIDTH-1 downto 0);
    vfpconfig_awprot          : out std_logic_vector(2 downto 0);
    vfpconfig_awvalid         : out std_logic;
    vfpconfig_awready         : in std_logic;
    vfpconfig_wdata           : out std_logic_vector(C_vfpConfig_DATA_WIDTH-1 downto 0);
    vfpconfig_wstrb           : out std_logic_vector((C_vfpConfig_DATA_WIDTH/8)-1 downto 0);
    vfpconfig_wvalid          : out std_logic;
    vfpconfig_wready          : in std_logic;
    vfpconfig_bresp           : in std_logic_vector(1 downto 0);
    vfpconfig_bvalid          : in std_logic;
    vfpconfig_bready          : out std_logic;
    vfpconfig_araddr          : out std_logic_vector(C_vfpconfig_ADDR_WIDTH-1 downto 0);
    vfpconfig_arprot          : out std_logic_vector(2 downto 0);
    vfpconfig_arvalid         : out std_logic;
    vfpconfig_arready         : in std_logic;
    vfpconfig_rdata           : in std_logic_vector(C_vfpConfig_DATA_WIDTH-1 downto 0);
    vfpconfig_rresp           : in std_logic_vector(1 downto 0);
    vfpconfig_rvalid          : in std_logic;
    vfpconfig_rready          : out std_logic);
end dut_configAxis;
architecture arch_imp of dut_configAxis is
    -------------------------------------------------------------------------  
    constant configRegister1                      : integer := 0;
    constant configRegister2                      : integer := 4;
    constant configRegister3                      : integer := 8;
    constant aBusSelect                           : integer := 12;
    constant configRegister5                      : integer := 16;
    constant videoChannel                         : integer := 20;
    constant dChannel                             : integer := 24;
    constant configRegister8                      : integer := 28;
    constant configRegister9                      : integer := 32;
    constant configRegister10                     : integer := 36;
    constant configRegister11                     : integer := 40;
    constant configRegister12                     : integer := 44;
    constant configRegister13                     : integer := 48;
    constant configRegister14                     : integer := 52;
    constant configRegister15                     : integer := 56;
    constant configRegister16                     : integer := 60;
    constant configRegister17                     : integer := 64;
    constant configRegister18                     : integer := 68;
    constant configRegister19                     : integer := 72;
    constant configRegister20                     : integer := 76;
    constant configRegister21                     : integer := 80;
    constant configRegister22                     : integer := 84;
    constant configRegister23                     : integer := 88;
    constant configRegister24                     : integer := 92;
    constant configRegister25                     : integer := 96;
    constant configRegister26                     : integer := 100;
    constant configRegister27                     : integer := 104;
    constant configRegister28                     : integer := 108;
    constant configRegister29                     : integer := 112;
    constant configRegister30                     : integer := 116;
    constant configRegister31                     : integer := 120;
    constant configRegister32                     : integer := 124;
	constant configRegister33	                  : integer := 128;
	constant configRegister34	                  : integer := 132;
	constant configRegister35	                  : integer := 136;
	constant configRegister36	                  : integer := 140;
	constant configRegister37	                  : integer := 144;
	constant configRegister38	                  : integer := 148;
	constant configRegister39	                  : integer := 152;
	constant configRegister40	                  : integer := 156;
	constant configRegister41	                  : integer := 160;
	constant configRegister42	                  : integer := 164;
	constant configRegister43	                  : integer := 168;
	constant configRegister44	                  : integer := 172;
	constant configRegister45	                  : integer := 176;
	constant configRegister46	                  : integer := 180;
	constant configRegister47	                  : integer := 184;
	constant configRegister48	                  : integer := 188;
	constant configRegister49	                  : integer := 192;
	constant configRegister50	                  : integer := 196;
	constant configRegister51	                  : integer := 200;
	constant configRegister52	                  : integer := 204;
	constant configRegister53	                  : integer := 208;
	constant configRegister54	                  : integer := 212;
	constant configRegister55	                  : integer := 216;
	constant configRegister56	                  : integer := 220;
	constant configRegister57	                  : integer := 224;
	constant configRegister58	                  : integer := 228;
	constant configRegister59	                  : integer := 232;
	constant configRegister60	                  : integer := 236;
	constant configRegister61	                  : integer := 240;
	constant configRegister62	                  : integer := 244;
	constant configRegister63	                  : integer := 248;
	constant configRegister64	                  : integer := 252;
    -------------------------------------------------------------------------
    procedure maxi_write(
    constant Mawaddr    : integer;
    constant Mwdata     : integer;
    signal Maxi_awaddr  : out std_logic_vector(7 downto 0);
    signal Maxi_wdata   : out std_logic_vector(31 downto 0);
    signal Maxi_awvalid : out std_logic;
    signal Maxi_wvalid  : out std_logic;
    signal Maxi_awready : in std_logic;--address ready
    signal Maxi_wready  : in std_logic;--data ready
    signal Maxi_bready  : out std_logic;
    signal Maxi_bvalid  : in std_logic) is
    begin
        Maxi_awaddr  <= std_logic_vector(to_unsigned(Mawaddr, 8));
        Maxi_wdata   <= std_logic_vector(to_unsigned(Mwdata, Maxi_wdata'length));
        Maxi_awvalid <= '1';
        Maxi_wvalid  <= '1';
        wait until (Maxi_awready and Maxi_wready) = '1';
        Maxi_bready  <='1';
        wait until Maxi_bvalid = '1';  -- Write result valid
        Maxi_awvalid <= '0';
        Maxi_wvalid <= '0';
        Maxi_bready <= '1';
        wait until Maxi_bvalid = '0';-- All finished
        Maxi_bready <= '0';
    end procedure;
    -------------------------------------------------------------------------
    procedure maxi_read(
        constant araddr    : integer;
        signal axi_araddr  : out std_logic_vector(7 downto 0);
        signal axi_arready : in std_logic;
        signal axi_arvalid : out std_logic;
        signal axi_rready  : out std_logic;
        signal axi_rvalid  : in std_logic) is
        begin
            axi_araddr  <= std_logic_vector(to_unsigned(araddr, axi_araddr'length));
            axi_arvalid <= '1';
            axi_rready  <= '1';
            wait until axi_arready = '1';
            wait until axi_rvalid  = '1';
            axi_arvalid <= '0';
            axi_rready  <= '0';
    end procedure;
    -------------------------------------------------------------------------
    begin
    clk_gen(vfpconfig_aclk, aclk_freq);
    process begin
        vfpconfig_aresetn  <= '0';
    wait for 100 ns;
        vfpconfig_aresetn  <= '1';
    wait;
    end process;
    process begin
    vfpconfig_wstrb <=X"F";
    -------------------------------------------------------------------------------------------
    -- maxi_write(configRegister1,8,vfpconfig_awaddr,vfpconfig_wdata,vfpconfig_awvalid,vfpconfig_wvalid,vfpconfig_awready,vfpconfig_wready,vfpconfig_bready,vfpconfig_bvalid);
    -- maxi_write(configRegister2,16,vfpconfig_awaddr,vfpconfig_wdata,vfpconfig_awvalid,vfpconfig_wvalid,vfpconfig_awready,vfpconfig_wready,vfpconfig_bready,vfpconfig_bvalid);
    -- maxi_write(configRegister3,32,vfpconfig_awaddr,vfpconfig_wdata,vfpconfig_awvalid,vfpconfig_wvalid,vfpconfig_awready,vfpconfig_wready,vfpconfig_bready,vfpconfig_bvalid);
    -- maxi_write(aBusSelect,64,vfpconfig_awaddr,vfpconfig_wdata,vfpconfig_awvalid,vfpconfig_wvalid,vfpconfig_awready,vfpconfig_wready,vfpconfig_bready,vfpconfig_bvalid); 
    -- maxi_write(configRegister5,98,vfpconfig_awaddr,vfpconfig_wdata,vfpconfig_awvalid,vfpconfig_wvalid,vfpconfig_awready,vfpconfig_wready,vfpconfig_bready,vfpconfig_bvalid);
    -- maxi_write(videoChannel,3,vfpconfig_awaddr,vfpconfig_wdata,vfpconfig_awvalid,vfpconfig_wvalid,vfpconfig_awready,vfpconfig_wready,vfpconfig_bready,vfpconfig_bvalid);
    -- maxi_write(dChannel,1,vfpconfig_awaddr,vfpconfig_wdata,vfpconfig_awvalid,vfpconfig_wvalid,vfpconfig_awready,vfpconfig_wready,vfpconfig_bready,vfpconfig_bvalid);
    -- maxi_write(configRegister8,0,vfpconfig_awaddr,vfpconfig_wdata,vfpconfig_awvalid,vfpconfig_wvalid,vfpconfig_awready,vfpconfig_wready,vfpconfig_bready,vfpconfig_bvalid); 
    -- maxi_write(configRegister9,5,vfpconfig_awaddr,vfpconfig_wdata,vfpconfig_awvalid,vfpconfig_wvalid,vfpconfig_awready,vfpconfig_wready,vfpconfig_bready,vfpconfig_bvalid);
    -- maxi_write(configRegister10,16,vfpconfig_awaddr,vfpconfig_wdata,vfpconfig_awvalid,vfpconfig_wvalid,vfpconfig_awready,vfpconfig_wready,vfpconfig_bready,vfpconfig_bvalid);
    -- maxi_write(configRegister11,32,vfpconfig_awaddr,vfpconfig_wdata,vfpconfig_awvalid,vfpconfig_wvalid,vfpconfig_awready,vfpconfig_wready,vfpconfig_bready,vfpconfig_bvalid);
    -- maxi_write(configRegister12,64,vfpconfig_awaddr,vfpconfig_wdata,vfpconfig_awvalid,vfpconfig_wvalid,vfpconfig_awready,vfpconfig_wready,vfpconfig_bready,vfpconfig_bvalid); 
    -- maxi_write(configRegister13,8,vfpconfig_awaddr,vfpconfig_wdata,vfpconfig_awvalid,vfpconfig_wvalid,vfpconfig_awready,vfpconfig_wready,vfpconfig_bready,vfpconfig_bvalid);
    -- maxi_write(configRegister14,16,vfpconfig_awaddr,vfpconfig_wdata,vfpconfig_awvalid,vfpconfig_wvalid,vfpconfig_awready,vfpconfig_wready,vfpconfig_bready,vfpconfig_bvalid);
    -- maxi_write(configRegister15,32,vfpconfig_awaddr,vfpconfig_wdata,vfpconfig_awvalid,vfpconfig_wvalid,vfpconfig_awready,vfpconfig_wready,vfpconfig_bready,vfpconfig_bvalid);
    -- maxi_write(configRegister16,64,vfpconfig_awaddr,vfpconfig_wdata,vfpconfig_awvalid,vfpconfig_wvalid,vfpconfig_awready,vfpconfig_wready,vfpconfig_bready,vfpconfig_bvalid); 
    -- maxi_write(configRegister17,8,vfpconfig_awaddr,vfpconfig_wdata,vfpconfig_awvalid,vfpconfig_wvalid,vfpconfig_awready,vfpconfig_wready,vfpconfig_bready,vfpconfig_bvalid);
    -- maxi_write(configRegister18,16,vfpconfig_awaddr,vfpconfig_wdata,vfpconfig_awvalid,vfpconfig_wvalid,vfpconfig_awready,vfpconfig_wready,vfpconfig_bready,vfpconfig_bvalid);
    -- maxi_write(configRegister19,0,vfpconfig_awaddr,vfpconfig_wdata,vfpconfig_awvalid,vfpconfig_wvalid,vfpconfig_awready,vfpconfig_wready,vfpconfig_bready,vfpconfig_bvalid);
    -- maxi_write(configRegister20,127,vfpconfig_awaddr,vfpconfig_wdata,vfpconfig_awvalid,vfpconfig_wvalid,vfpconfig_awready,vfpconfig_wready,vfpconfig_bready,vfpconfig_bvalid); 
    -- maxi_write(configRegister21,7,vfpconfig_awaddr,vfpconfig_wdata,vfpconfig_awvalid,vfpconfig_wvalid,vfpconfig_awready,vfpconfig_wready,vfpconfig_bready,vfpconfig_bvalid);
    --pRegion.cpuWgridLock
    maxi_write(videoChannel,4,vfpconfig_awaddr,vfpconfig_wdata,vfpconfig_awvalid,vfpconfig_wvalid,vfpconfig_awready,vfpconfig_wready,vfpconfig_bready,vfpconfig_bvalid);
    maxi_write(dChannel,0,vfpconfig_awaddr,vfpconfig_wdata,vfpconfig_awvalid,vfpconfig_wvalid,vfpconfig_awready,vfpconfig_wready,vfpconfig_bready,vfpconfig_bvalid); 
    maxi_write(aBusSelect,3,vfpconfig_awaddr,vfpconfig_wdata,vfpconfig_awvalid,vfpconfig_wvalid,vfpconfig_awready,vfpconfig_wready,vfpconfig_bready,vfpconfig_bvalid); 
    maxi_write(configRegister31,0,vfpconfig_awaddr,vfpconfig_wdata,vfpconfig_awvalid,vfpconfig_wvalid,vfpconfig_awready,vfpconfig_wready,vfpconfig_bready,vfpconfig_bvalid); 
    maxi_write(configRegister35,1,vfpconfig_awaddr,vfpconfig_wdata,vfpconfig_awvalid,vfpconfig_wvalid,vfpconfig_awready,vfpconfig_wready,vfpconfig_bready,vfpconfig_bvalid); 
    maxi_write(configRegister8,1,vfpconfig_awaddr,vfpconfig_wdata,vfpconfig_awvalid,vfpconfig_wvalid,vfpconfig_awready,vfpconfig_wready,vfpconfig_bready,vfpconfig_bvalid); 
    maxi_write(configRegister40,1,vfpconfig_awaddr,vfpconfig_wdata,vfpconfig_awvalid,vfpconfig_wvalid,vfpconfig_awready,vfpconfig_wready,vfpconfig_bready,vfpconfig_bvalid); 
    maxi_write(configRegister40,0,vfpconfig_awaddr,vfpconfig_wdata,vfpconfig_awvalid,vfpconfig_wvalid,vfpconfig_awready,vfpconfig_wready,vfpconfig_bready,vfpconfig_bvalid); 
    maxi_write(configRegister32,10,vfpconfig_awaddr,vfpconfig_wdata,vfpconfig_awvalid,vfpconfig_wvalid,vfpconfig_awready,vfpconfig_wready,vfpconfig_bready,vfpconfig_bvalid); 
    wait for 500 us;
    maxi_write(configRegister37,0,vfpconfig_awaddr,vfpconfig_wdata,vfpconfig_awvalid,vfpconfig_wvalid,vfpconfig_awready,vfpconfig_wready,vfpconfig_bready,vfpconfig_bvalid);
    maxi_read(configRegister39, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    maxi_write(configRegister37,1,vfpconfig_awaddr,vfpconfig_wdata,vfpconfig_awvalid,vfpconfig_wvalid,vfpconfig_awready,vfpconfig_wready,vfpconfig_bready,vfpconfig_bvalid);
    maxi_read(configRegister39, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    maxi_write(configRegister37,2,vfpconfig_awaddr,vfpconfig_wdata,vfpconfig_awvalid,vfpconfig_wvalid,vfpconfig_awready,vfpconfig_wready,vfpconfig_bready,vfpconfig_bvalid);
    maxi_read(configRegister39, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    maxi_write(configRegister37,3,vfpconfig_awaddr,vfpconfig_wdata,vfpconfig_awvalid,vfpconfig_wvalid,vfpconfig_awready,vfpconfig_wready,vfpconfig_bready,vfpconfig_bvalid);
    maxi_read(configRegister39, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    maxi_write(configRegister37,4,vfpconfig_awaddr,vfpconfig_wdata,vfpconfig_awvalid,vfpconfig_wvalid,vfpconfig_awready,vfpconfig_wready,vfpconfig_bready,vfpconfig_bvalid);
    maxi_read(configRegister39, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_write(configRegister23,32,vfpconfig_awaddr,vfpconfig_wdata,vfpconfig_awvalid,vfpconfig_wvalid,vfpconfig_awready,vfpconfig_wready,vfpconfig_bready,vfpconfig_bvalid);
    -- maxi_write(configRegister24,64,vfpconfig_awaddr,vfpconfig_wdata,vfpconfig_awvalid,vfpconfig_wvalid,vfpconfig_awready,vfpconfig_wready,vfpconfig_bready,vfpconfig_bvalid); 
    -- maxi_write(configRegister25,8,vfpconfig_awaddr,vfpconfig_wdata,vfpconfig_awvalid,vfpconfig_wvalid,vfpconfig_awready,vfpconfig_wready,vfpconfig_bready,vfpconfig_bvalid);
    -- maxi_write(configRegister26,16,vfpconfig_awaddr,vfpconfig_wdata,vfpconfig_awvalid,vfpconfig_wvalid,vfpconfig_awready,vfpconfig_wready,vfpconfig_bready,vfpconfig_bvalid);
    -- maxi_write(configRegister27,32,vfpconfig_awaddr,vfpconfig_wdata,vfpconfig_awvalid,vfpconfig_wvalid,vfpconfig_awready,vfpconfig_wready,vfpconfig_bready,vfpconfig_bvalid);
    -- maxi_write(configRegister28,64,vfpconfig_awaddr,vfpconfig_wdata,vfpconfig_awvalid,vfpconfig_wvalid,vfpconfig_awready,vfpconfig_wready,vfpconfig_bready,vfpconfig_bvalid); 
    -- maxi_write(configRegister29,8,vfpconfig_awaddr,vfpconfig_wdata,vfpconfig_awvalid,vfpconfig_wvalid,vfpconfig_awready,vfpconfig_wready,vfpconfig_bready,vfpconfig_bvalid);
    -- maxi_write(configRegister30,16,vfpconfig_awaddr,vfpconfig_wdata,vfpconfig_awvalid,vfpconfig_wvalid,vfpconfig_awready,vfpconfig_wready,vfpconfig_bready,vfpconfig_bvalid);
    -- maxi_write(configRegister31,32,vfpconfig_awaddr,vfpconfig_wdata,vfpconfig_awvalid,vfpconfig_wvalid,vfpconfig_awready,vfpconfig_wready,vfpconfig_bready,vfpconfig_bvalid);
    -- maxi_write(configRegister32,64,vfpconfig_awaddr,vfpconfig_wdata,vfpconfig_awvalid,vfpconfig_wvalid,vfpconfig_awready,vfpconfig_wready,vfpconfig_bready,vfpconfig_bvalid);
    -------------------------------------------------------------------------------------------
    -- maxi_read(configRegister1, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister2, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister1, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister2, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister1, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister2, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister1, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister2, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister1, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister2, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister1, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister2, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister1, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister2, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister1, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister2, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister1, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister2, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister1, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister2, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister1, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister2, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister1, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister2, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister1, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister2, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister1, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister2, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister1, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister2, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister1, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister2, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister1, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister2, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister1, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister2, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister1, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister2, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister1, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister2, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister1, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister2, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister1, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister2, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister1, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister2, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister1, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister2, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister1, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister2, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister1, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister2, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister1, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister2, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister1, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister2, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister1, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister2, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister1, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister2, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister1, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister2, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister1, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister2, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister1, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister2, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister1, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister2, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister1, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister2, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister1, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister2, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister1, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister2, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister1, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister2, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister1, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister2, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister1, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister2, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister1, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister2, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister1, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister2, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister1, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister2, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister1, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister2, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister1, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister2, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister1, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister2, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister1, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister2, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister1, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister2, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister1, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister2, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister1, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister2, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister1, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister2, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister1, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister2, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister1, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister2, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister1, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister2, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister1, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister2, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister1, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister2, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister1, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister2, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister1, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister2, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister1, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister2, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister3, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(aBusSelect, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister5, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(videoChannel, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister7, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister8, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister9, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister10, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister11, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister12, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister13, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister14, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister15, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister16, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister17, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister18, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister19, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister20, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister21, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister22, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister23, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister24, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister25, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister26, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister27, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister28, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    -- maxi_read(configRegister29, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
     --maxi_read(configRegister30, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
     --maxi_read(configRegister31, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
     --maxi_read(configRegister32, vfpconfig_araddr, vfpconfig_arready, vfpconfig_arvalid, vfpconfig_rready, vfpconfig_rvalid);
    wait;
    end process;
end arch_imp;