// Class: img_seqr
typedef uvm_sequencer #(d5m_trans) img_seqr; 
//class img_seqr extends uvm_sequencer #(d5m_trans);
//
//    int id;
//    
//    `uvm_component_utils_begin(img_seqr)
//        `uvm_field_int(id, UVM_DEFAULT)
//    `uvm_component_utils_end
//    
//    // Function: new
//    function new (string name, uvm_component parent);
//        super.new(name, parent);
//    endfunction: new
//    
//endclass: img_seqr