-------------------------------------------------------------------------------
--
-- Filename    : d_valid.vhd
-- Create Date : 01162019 [01-16-2019]
-- Author      : Zakinder
--
-- Description:
-- This file instantiation
--
-------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.constants_package.all;
use work.vpf_records.all;
use work.ports_package.all;
entity d_valid is
generic (
    pixelDelay     : integer := 8);
port (
    clk            : in std_logic;
    iRgb           : in channel;
    oRgb           : out channel);
end d_valid;
architecture behavioral of d_valid is
signal rgbSyncValid    : std_logic_vector(56 downto 0)  := (others => '0');
signal rgbSyncEol      : std_logic_vector(56 downto 0)  := (others => '0');
signal rgbSyncSof      : std_logic_vector(56 downto 0)  := (others => '0');
signal rgbSyncEof      : std_logic_vector(56 downto 0)  := (others => '0');
begin
process (clk) begin
    if rising_edge(clk) then
        rgbSyncValid(0)  <= iRgb.valid;
        rgbSyncValid(1)  <= rgbSyncValid(0);
        rgbSyncValid(2)  <= rgbSyncValid(1);
        rgbSyncValid(3)  <= rgbSyncValid(2);
        rgbSyncValid(4)  <= rgbSyncValid(3);
        rgbSyncValid(5)  <= rgbSyncValid(4);
        rgbSyncValid(6)  <= rgbSyncValid(5);
        rgbSyncValid(7)  <= rgbSyncValid(6);
        rgbSyncValid(8)  <= rgbSyncValid(7);
        rgbSyncValid(9)  <= rgbSyncValid(8);
        rgbSyncValid(10) <= rgbSyncValid(9);
        rgbSyncValid(11) <= rgbSyncValid(10);
        rgbSyncValid(12) <= rgbSyncValid(11);
        rgbSyncValid(13) <= rgbSyncValid(12);
        rgbSyncValid(14) <= rgbSyncValid(13);
        rgbSyncValid(15) <= rgbSyncValid(14);
        rgbSyncValid(16) <= rgbSyncValid(15);
        rgbSyncValid(17) <= rgbSyncValid(16);
        rgbSyncValid(18) <= rgbSyncValid(17);
        rgbSyncValid(19) <= rgbSyncValid(18);
        rgbSyncValid(20) <= rgbSyncValid(19);
        rgbSyncValid(21) <= rgbSyncValid(20);
        rgbSyncValid(22) <= rgbSyncValid(21);
        rgbSyncValid(23) <= rgbSyncValid(22);
        rgbSyncValid(24) <= rgbSyncValid(23);
        rgbSyncValid(25) <= rgbSyncValid(24);
        rgbSyncValid(26) <= rgbSyncValid(25);
        rgbSyncValid(27) <= rgbSyncValid(26);
        rgbSyncValid(28) <= rgbSyncValid(27);
        rgbSyncValid(29) <= rgbSyncValid(28);
        rgbSyncValid(30) <= rgbSyncValid(29);
        rgbSyncValid(31) <= rgbSyncValid(30);
        rgbSyncValid(32) <= rgbSyncValid(31);
        rgbSyncValid(33) <= rgbSyncValid(32);
        rgbSyncValid(34) <= rgbSyncValid(33);
        rgbSyncValid(35) <= rgbSyncValid(34);
        rgbSyncValid(36) <= rgbSyncValid(35);
        rgbSyncValid(37) <= rgbSyncValid(36);
        rgbSyncValid(38) <= rgbSyncValid(37);
        rgbSyncValid(39) <= rgbSyncValid(38);
        rgbSyncValid(40) <= rgbSyncValid(39);
        rgbSyncValid(41) <= rgbSyncValid(40);
        rgbSyncValid(42) <= rgbSyncValid(41);
        rgbSyncValid(43) <= rgbSyncValid(42);
        rgbSyncValid(44) <= rgbSyncValid(43);
        rgbSyncValid(45) <= rgbSyncValid(44);
        rgbSyncValid(46) <= rgbSyncValid(45);
        rgbSyncValid(47) <= rgbSyncValid(46);
        rgbSyncValid(48) <= rgbSyncValid(47);
        rgbSyncValid(49) <= rgbSyncValid(48);
        rgbSyncValid(50) <= rgbSyncValid(49);
        rgbSyncValid(51) <= rgbSyncValid(50);
        rgbSyncValid(52) <= rgbSyncValid(51);
        rgbSyncValid(53) <= rgbSyncValid(52);
        rgbSyncValid(54) <= rgbSyncValid(53);
        rgbSyncValid(55) <= rgbSyncValid(54);
        rgbSyncValid(56) <= rgbSyncValid(55);
    end if;
end process;
process (clk) begin
    if rising_edge(clk) then
        rgbSyncEol(0)  <= iRgb.eol;
        rgbSyncEol(1)  <= rgbSyncEol(0);
        rgbSyncEol(2)  <= rgbSyncEol(1);
        rgbSyncEol(3)  <= rgbSyncEol(2);
        rgbSyncEol(4)  <= rgbSyncEol(3);
        rgbSyncEol(5)  <= rgbSyncEol(4);
        rgbSyncEol(6)  <= rgbSyncEol(5);
        rgbSyncEol(7)  <= rgbSyncEol(6);
        rgbSyncEol(8)  <= rgbSyncEol(7);
        rgbSyncEol(9)  <= rgbSyncEol(8);
        rgbSyncEol(10) <= rgbSyncEol(9);
        rgbSyncEol(11) <= rgbSyncEol(10);
        rgbSyncEol(12) <= rgbSyncEol(11);
        rgbSyncEol(13) <= rgbSyncEol(12);
        rgbSyncEol(14) <= rgbSyncEol(13);
        rgbSyncEol(15) <= rgbSyncEol(14);
        rgbSyncEol(16) <= rgbSyncEol(15);
        rgbSyncEol(17) <= rgbSyncEol(16);
        rgbSyncEol(18) <= rgbSyncEol(17);
        rgbSyncEol(19) <= rgbSyncEol(18);
        rgbSyncEol(20) <= rgbSyncEol(19);
        rgbSyncEol(21) <= rgbSyncEol(20);
        rgbSyncEol(22) <= rgbSyncEol(21);
        rgbSyncEol(23) <= rgbSyncEol(22);
        rgbSyncEol(24) <= rgbSyncEol(23);
        rgbSyncEol(25) <= rgbSyncEol(24);
        rgbSyncEol(26) <= rgbSyncEol(25);
        rgbSyncEol(27) <= rgbSyncEol(26);
        rgbSyncEol(28) <= rgbSyncEol(27);
        rgbSyncEol(29) <= rgbSyncEol(28);
        rgbSyncEol(30) <= rgbSyncEol(29);
        rgbSyncEol(31) <= rgbSyncEol(30);
        rgbSyncEol(32) <= rgbSyncEol(31);
        rgbSyncEol(33) <= rgbSyncEol(32);
        rgbSyncEol(34) <= rgbSyncEol(33);
        rgbSyncEol(35) <= rgbSyncEol(34);
        rgbSyncEol(36) <= rgbSyncEol(35);
        rgbSyncEol(37) <= rgbSyncEol(36);
        rgbSyncEol(38) <= rgbSyncEol(37);
        rgbSyncEol(39) <= rgbSyncEol(38);
        rgbSyncEol(40) <= rgbSyncEol(39);
        rgbSyncEol(41) <= rgbSyncEol(40);
        rgbSyncEol(42) <= rgbSyncEol(41);
        rgbSyncEol(43) <= rgbSyncEol(42);
        rgbSyncEol(44) <= rgbSyncEol(43);
        rgbSyncEol(45) <= rgbSyncEol(44);
        rgbSyncEol(46) <= rgbSyncEol(45);
        rgbSyncEol(47) <= rgbSyncEol(46);
        rgbSyncEol(48) <= rgbSyncEol(47);
        rgbSyncEol(49) <= rgbSyncEol(48);
        rgbSyncEol(50) <= rgbSyncEol(49);
        rgbSyncEol(51) <= rgbSyncEol(50);
        rgbSyncEol(52) <= rgbSyncEol(51);
        rgbSyncEol(53) <= rgbSyncEol(52);
        rgbSyncEol(54) <= rgbSyncEol(53);
        rgbSyncEol(55) <= rgbSyncEol(54);
        rgbSyncEol(56) <= rgbSyncEol(55);
    end if;
end process;
process (clk) begin
    if rising_edge(clk) then
        rgbSyncSof(0)  <= iRgb.sof;
        rgbSyncSof(1)  <= rgbSyncSof(0);
        rgbSyncSof(2)  <= rgbSyncSof(1);
        rgbSyncSof(3)  <= rgbSyncSof(2);
        rgbSyncSof(4)  <= rgbSyncSof(3);
        rgbSyncSof(5)  <= rgbSyncSof(4);
        rgbSyncSof(6)  <= rgbSyncSof(5);
        rgbSyncSof(7)  <= rgbSyncSof(6);
        rgbSyncSof(8)  <= rgbSyncSof(7);
        rgbSyncSof(9)  <= rgbSyncSof(8);
        rgbSyncSof(10) <= rgbSyncSof(9);
        rgbSyncSof(11) <= rgbSyncSof(10);
        rgbSyncSof(12) <= rgbSyncSof(11);
        rgbSyncSof(13) <= rgbSyncSof(12);
        rgbSyncSof(14) <= rgbSyncSof(13);
        rgbSyncSof(15) <= rgbSyncSof(14);
        rgbSyncSof(16) <= rgbSyncSof(15);
        rgbSyncSof(17) <= rgbSyncSof(16);
        rgbSyncSof(18) <= rgbSyncSof(17);
        rgbSyncSof(19) <= rgbSyncSof(18);
        rgbSyncSof(20) <= rgbSyncSof(19);
        rgbSyncSof(21) <= rgbSyncSof(20);
        rgbSyncSof(22) <= rgbSyncSof(21);
        rgbSyncSof(23) <= rgbSyncSof(22);
        rgbSyncSof(24) <= rgbSyncSof(23);
        rgbSyncSof(25) <= rgbSyncSof(24);
        rgbSyncSof(26) <= rgbSyncSof(25);
        rgbSyncSof(27) <= rgbSyncSof(26);
        rgbSyncSof(28) <= rgbSyncSof(27);
        rgbSyncSof(29) <= rgbSyncSof(28);
        rgbSyncSof(30) <= rgbSyncSof(29);
        rgbSyncSof(31) <= rgbSyncSof(30);
        rgbSyncSof(32) <= rgbSyncSof(31);
        rgbSyncSof(33) <= rgbSyncSof(32);
        rgbSyncSof(34) <= rgbSyncSof(33);
        rgbSyncSof(35) <= rgbSyncSof(34);
        rgbSyncSof(36) <= rgbSyncSof(35);
        rgbSyncSof(37) <= rgbSyncSof(36);
        rgbSyncSof(38) <= rgbSyncSof(37);
        rgbSyncSof(39) <= rgbSyncSof(38);
        rgbSyncSof(40) <= rgbSyncSof(39);
        rgbSyncSof(41) <= rgbSyncSof(40);
        rgbSyncSof(42) <= rgbSyncSof(41);
        rgbSyncSof(43) <= rgbSyncSof(42);
        rgbSyncSof(44) <= rgbSyncSof(43);
        rgbSyncSof(45) <= rgbSyncSof(44);
        rgbSyncSof(46) <= rgbSyncSof(45);
        rgbSyncSof(47) <= rgbSyncSof(46);
        rgbSyncSof(48) <= rgbSyncSof(47);
        rgbSyncSof(49) <= rgbSyncSof(48);
        rgbSyncSof(50) <= rgbSyncSof(49);
        rgbSyncSof(51) <= rgbSyncSof(50);
        rgbSyncSof(52) <= rgbSyncSof(51);
        rgbSyncSof(53) <= rgbSyncSof(52);
        rgbSyncSof(54) <= rgbSyncSof(53);
        rgbSyncSof(55) <= rgbSyncSof(54);
        rgbSyncSof(56) <= rgbSyncSof(55);
    end if;
end process;
process (clk) begin
    if rising_edge(clk) then
        rgbSyncEof(0)  <= iRgb.eof;
        rgbSyncEof(1)  <= rgbSyncEof(0);
        rgbSyncEof(2)  <= rgbSyncEof(1);
        rgbSyncEof(3)  <= rgbSyncEof(2);
        rgbSyncEof(4)  <= rgbSyncEof(3);
        rgbSyncEof(5)  <= rgbSyncEof(4);
        rgbSyncEof(6)  <= rgbSyncEof(5);
        rgbSyncEof(7)  <= rgbSyncEof(6);
        rgbSyncEof(8)  <= rgbSyncEof(7);
        rgbSyncEof(9)  <= rgbSyncEof(8);
        rgbSyncEof(10) <= rgbSyncEof(9);
        rgbSyncEof(11) <= rgbSyncEof(10);
        rgbSyncEof(12) <= rgbSyncEof(11);
        rgbSyncEof(13) <= rgbSyncEof(12);
        rgbSyncEof(14) <= rgbSyncEof(13);
        rgbSyncEof(15) <= rgbSyncEof(14);
        rgbSyncEof(16) <= rgbSyncEof(15);
        rgbSyncEof(17) <= rgbSyncEof(16);
        rgbSyncEof(18) <= rgbSyncEof(17);
        rgbSyncEof(19) <= rgbSyncEof(18);
        rgbSyncEof(20) <= rgbSyncEof(19);
        rgbSyncEof(21) <= rgbSyncEof(20);
        rgbSyncEof(22) <= rgbSyncEof(21);
        rgbSyncEof(23) <= rgbSyncEof(22);
        rgbSyncEof(24) <= rgbSyncEof(23);
        rgbSyncEof(25) <= rgbSyncEof(24);
        rgbSyncEof(26) <= rgbSyncEof(25);
        rgbSyncEof(27) <= rgbSyncEof(26);
        rgbSyncEof(28) <= rgbSyncEof(27);
        rgbSyncEof(29) <= rgbSyncEof(28);
        rgbSyncEof(30) <= rgbSyncEof(29);
        rgbSyncEof(31) <= rgbSyncEof(30);
        rgbSyncEof(32) <= rgbSyncEof(31);
        rgbSyncEof(33) <= rgbSyncEof(32);
        rgbSyncEof(34) <= rgbSyncEof(33);
        rgbSyncEof(35) <= rgbSyncEof(34);
        rgbSyncEof(36) <= rgbSyncEof(35);
        rgbSyncEof(37) <= rgbSyncEof(36);
        rgbSyncEof(38) <= rgbSyncEof(37);
        rgbSyncEof(39) <= rgbSyncEof(38);
        rgbSyncEof(40) <= rgbSyncEof(39);
        rgbSyncEof(41) <= rgbSyncEof(40);
        rgbSyncEof(42) <= rgbSyncEof(41);
        rgbSyncEof(43) <= rgbSyncEof(42);
        rgbSyncEof(44) <= rgbSyncEof(43);
        rgbSyncEof(45) <= rgbSyncEof(44);
        rgbSyncEof(46) <= rgbSyncEof(45);
        rgbSyncEof(47) <= rgbSyncEof(46);
        rgbSyncEof(48) <= rgbSyncEof(47);
        rgbSyncEof(49) <= rgbSyncEof(48);
        rgbSyncEof(50) <= rgbSyncEof(49);
        rgbSyncEof(51) <= rgbSyncEof(50);
        rgbSyncEof(52) <= rgbSyncEof(51);
        rgbSyncEof(53) <= rgbSyncEof(52);
        rgbSyncEof(54) <= rgbSyncEof(53);
        rgbSyncEof(55) <= rgbSyncEof(54);
        rgbSyncEof(56) <= rgbSyncEof(55);
    end if;
end process;
    oRgb.red      <= iRgb.red;
    oRgb.green    <= iRgb.green;
    oRgb.blue     <= iRgb.blue;
    oRgb.valid    <= rgbSyncValid(pixelDelay);
    oRgb.eol      <= rgbSyncEol(pixelDelay);
    oRgb.sof      <= rgbSyncSof(pixelDelay);
    oRgb.eof      <= rgbSyncEof(pixelDelay);
end behavioral;