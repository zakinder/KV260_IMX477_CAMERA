-------------------------------------------------------------------------------
--
-- Filename    : rgb_range.vhd
-- Create Date : 02092019 [02-17-2019]
-- Author      : Zakinder
--
-- Description:
-- This file instantiation axi4 components.
--
-------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.constants_package.all;
use work.vpf_records.all;
use work.ports_package.all;
entity rgb_range is
generic (
    i_data_width      : integer := 8);
port (
    clk            : in  std_logic;
    reset          : in  std_logic;
    gain           : in  natural;
    iRgb           : in channel;
    oRgb           : out channel);
end rgb_range;
architecture Behavioral of rgb_range is
    signal i1Rgb       : intChannel;
    signal i2Rgb       : intChannel;
    signal i3Rgb       : intChannel;
    signal rgbSyncEol  : std_logic;
    signal rgbSyncSof  : std_logic;
    signal rgbSyncEof  : std_logic;
    --constant gain      : natural := 0;
    
begin

process (clk)begin
    if rising_edge(clk) then
        rgbSyncEol   <= iRgb.eol;
        rgbSyncSof   <= iRgb.sof;
        rgbSyncEof   <= iRgb.eof;
    end if;
end process;


process (clk,reset)begin
    if (reset = lo) then
        i1Rgb.red    <= zero;
        i1Rgb.green  <= zero;
        i1Rgb.blue   <= zero;
    elsif rising_edge(clk) then
        i1Rgb.red    <= to_integer(unsigned(iRgb.red));
        i1Rgb.green  <= to_integer(unsigned(iRgb.green));
        i1Rgb.blue   <= to_integer(unsigned(iRgb.blue));
        i1Rgb.valid  <= iRgb.valid;
        i2Rgb.valid  <= i1Rgb.valid;
        i3Rgb        <= i2Rgb;
    end if;
end process;
---------------------------------------------------------------------------------
-- i2Rgb.valid must be 2nd condition else valid value
---------------------------------------------------------------------------------
process (clk) begin
    if rising_edge(clk) then
      if (i1Rgb.red   >= 0 and     i1Rgb.red <= 9)               then  i2Rgb.red <= 7;
      elsif (i1Rgb.red   >= 10 and    i1Rgb.red <= (19))         then  i2Rgb.red <= 17;
      elsif (i1Rgb.red   >= 20 and    i1Rgb.red <= (29))         then  i2Rgb.red <= 27;
      elsif (i1Rgb.red   >= 30 and    i1Rgb.red <= (39+gain))    then  i2Rgb.red <= 37;
      elsif (i1Rgb.red   >= 40 and    i1Rgb.red <= (49+gain))    then  i2Rgb.red <= 47;
      elsif (i1Rgb.red   >= 50 and    i1Rgb.red <= (59+gain))    then  i2Rgb.red <= 57;
      elsif (i1Rgb.red   >= 60 and    i1Rgb.red <= (69+gain))    then  i2Rgb.red <= 67;
      elsif (i1Rgb.red   >= 70 and    i1Rgb.red <= (79+gain))    then  i2Rgb.red <= 77;
      elsif (i1Rgb.red   >= 80 and    i1Rgb.red <= (89+gain))    then  i2Rgb.red <= 87;
      elsif (i1Rgb.red   >= 90 and    i1Rgb.red <= (99+gain))    then  i2Rgb.red <= 97;
      elsif (i1Rgb.red   >= 100 and   i1Rgb.red <= (109+gain))   then  i2Rgb.red <= 107;
      elsif (i1Rgb.red   >= 110 and   i1Rgb.red <= (119+gain))   then  i2Rgb.red <= 117;
      elsif (i1Rgb.red   >= 120 and   i1Rgb.red <= (129+gain))   then  i2Rgb.red <= 127;
      elsif (i1Rgb.red   >= 130 and   i1Rgb.red <= (139+gain))   then  i2Rgb.red <= 137;
      elsif (i1Rgb.red   >= 140 and   i1Rgb.red <= (149+gain))   then  i2Rgb.red <= 147;
      elsif (i1Rgb.red   >= 150 and   i1Rgb.red <= (159+gain))   then  i2Rgb.red <= 157;
      elsif (i1Rgb.red   >= 160 and   i1Rgb.red <= (169+gain))   then  i2Rgb.red <= 167;
      elsif (i1Rgb.red   >= 170 and   i1Rgb.red <= (179+gain))   then  i2Rgb.red <= 177;
      elsif (i1Rgb.red   >= 180 and   i1Rgb.red <= (189+gain))   then  i2Rgb.red <= 187;
      elsif (i1Rgb.red   >= 190 and   i1Rgb.red <= (199+gain))   then  i2Rgb.red <= 197;
      elsif (i1Rgb.red   >= 200 and   i1Rgb.red <= (209+gain))   then  i2Rgb.red <= 207;
      elsif (i1Rgb.red   >= 210 and   i1Rgb.red <= (219+gain))   then  i2Rgb.red <= 217;
      elsif (i1Rgb.red   >= 220 and   i1Rgb.red <= (229+gain))   then  i2Rgb.red <= 227;
      elsif (i1Rgb.red   >= 230 and   i1Rgb.red <= (239+gain))   then  i2Rgb.red <= 237;
      elsif (i1Rgb.red   >= 240 and   i1Rgb.red <= (249+gain))   then  i2Rgb.red <= 247;
      elsif (i1Rgb.red   >= 250 and   i1Rgb.red <= (259+gain))   then  i2Rgb.red <= 257;
      elsif (i1Rgb.red   >= 260 and   i1Rgb.red <= (269+gain))   then  i2Rgb.red <= 267;
      elsif (i1Rgb.red   >= 270 and   i1Rgb.red <= (279+gain))   then  i2Rgb.red <= 277;
      elsif (i1Rgb.red   >= 280 and   i1Rgb.red <= (289+gain))   then  i2Rgb.red <= 287;
      elsif (i1Rgb.red   >= 290 and   i1Rgb.red <= (299+gain))   then  i2Rgb.red <= 297;
      elsif (i1Rgb.red   >= 300 and   i1Rgb.red <= (309+gain))   then  i2Rgb.red <= 307;
      elsif (i1Rgb.red   >= 310 and   i1Rgb.red <= (319+gain))   then  i2Rgb.red <= 317;
      elsif (i1Rgb.red   >= 320 and   i1Rgb.red <= (329+gain))   then  i2Rgb.red <= 327;
      elsif (i1Rgb.red   >= 330 and   i1Rgb.red <= (339+gain))   then  i2Rgb.red <= 337;
      elsif (i1Rgb.red   >= 340 and   i1Rgb.red <= (349+gain))   then  i2Rgb.red <= 347;
      elsif (i1Rgb.red   >= 350 and   i1Rgb.red <= (359+gain))   then  i2Rgb.red <= 357;
      elsif (i1Rgb.red   >= 360 and   i1Rgb.red <= (369+gain))   then  i2Rgb.red <= 367;
      elsif (i1Rgb.red   >= 370 and   i1Rgb.red <= (379+gain))   then  i2Rgb.red <= 377;
      elsif (i1Rgb.red   >= 380 and   i1Rgb.red <= (389+gain))   then  i2Rgb.red <= 387;
      elsif (i1Rgb.red   >= 390 and   i1Rgb.red <= (399+gain))   then  i2Rgb.red <= 397;
      elsif (i1Rgb.red   >= 400 and   i1Rgb.red <= (409+gain))   then  i2Rgb.red <= 407;
      elsif (i1Rgb.red   >= 400 and   i1Rgb.red <= (409+gain))   then  i2Rgb.red <= 407;
      elsif (i1Rgb.red   >= 410 and   i1Rgb.red <= (419+gain))   then  i2Rgb.red <= 417;
      elsif (i1Rgb.red   >= 420 and   i1Rgb.red <= (429+gain))   then  i2Rgb.red <= 427;
      elsif (i1Rgb.red   >= 430 and   i1Rgb.red <= (439+gain))   then  i2Rgb.red <= 437;
      elsif (i1Rgb.red   >= 440 and   i1Rgb.red <= (449+gain))   then  i2Rgb.red <= 447;
      elsif (i1Rgb.red   >= 450 and   i1Rgb.red <= (459+gain))   then  i2Rgb.red <= 457;
      elsif (i1Rgb.red   >= 460 and   i1Rgb.red <= (469+gain))   then  i2Rgb.red <= 467;
      elsif (i1Rgb.red   >= 470 and   i1Rgb.red <= (479+gain))   then  i2Rgb.red <= 477;
      elsif (i1Rgb.red   >= 480 and   i1Rgb.red <= (489+gain))   then  i2Rgb.red <= 487;
      elsif (i1Rgb.red   >= 490 and   i1Rgb.red <= (499+gain))   then  i2Rgb.red <= 497;
      elsif (i1Rgb.red   >= 500 and   i1Rgb.red <= (509+gain))   then  i2Rgb.red <= 507;
      elsif (i1Rgb.red   >= 510 and   i1Rgb.red <= (519+gain))   then  i2Rgb.red <= 517;
      elsif (i1Rgb.red   >= 520 and   i1Rgb.red <= (529+gain))   then  i2Rgb.red <= 527;
      elsif (i1Rgb.red   >= 530 and   i1Rgb.red <= (539+gain))   then  i2Rgb.red <= 537;
      elsif (i1Rgb.red   >= 540 and   i1Rgb.red <= (549+gain))   then  i2Rgb.red <= 547;
      elsif (i1Rgb.red   >= 550 and   i1Rgb.red <= (559+gain))   then  i2Rgb.red <= 557;
      elsif (i1Rgb.red   >= 560 and   i1Rgb.red <= (569+gain))   then  i2Rgb.red <= 567;
      elsif (i1Rgb.red   >= 570 and   i1Rgb.red <= (579+gain))   then  i2Rgb.red <= 577;
      elsif (i1Rgb.red   >= 580 and   i1Rgb.red <= (589+gain))   then  i2Rgb.red <= 587;
      elsif (i1Rgb.red   >= 590 and   i1Rgb.red <= (599+gain))   then  i2Rgb.red <= 597;
      elsif (i1Rgb.red   >= 600 and   i1Rgb.red <= (609+gain))   then  i2Rgb.red <= 607;
      elsif (i1Rgb.red   >= 610 and   i1Rgb.red <= (619+gain))   then  i2Rgb.red <= 617;
      elsif (i1Rgb.red   >= 620 and   i1Rgb.red <= (629+gain))   then  i2Rgb.red <= 627;
      elsif (i1Rgb.red   >= 630 and   i1Rgb.red <= (639+gain))   then  i2Rgb.red <= 637;
      elsif (i1Rgb.red   >= 640 and   i1Rgb.red <= (649+gain))   then  i2Rgb.red <= 647;
      elsif (i1Rgb.red   >= 650 and   i1Rgb.red <= (659+gain))   then  i2Rgb.red <= 657;
      elsif (i1Rgb.red   >= 660 and   i1Rgb.red <= (669+gain))   then  i2Rgb.red <= 667;
      elsif (i1Rgb.red   >= 670 and   i1Rgb.red <= (679+gain))   then  i2Rgb.red <= 677;
      elsif (i1Rgb.red   >= 680 and   i1Rgb.red <= (689+gain))   then  i2Rgb.red <= 687;
      elsif (i1Rgb.red   >= 690 and   i1Rgb.red <= (699+gain))   then  i2Rgb.red <= 697;
      elsif (i1Rgb.red   >= 700 and   i1Rgb.red <= (709+gain))   then  i2Rgb.red <= 707;
      elsif (i1Rgb.red   >= 710 and   i1Rgb.red <= (719+gain))   then  i2Rgb.red <= 717;
      elsif (i1Rgb.red   >= 720 and   i1Rgb.red <= (729+gain))   then  i2Rgb.red <= 727;
      elsif (i1Rgb.red   >= 730 and   i1Rgb.red <= (739+gain))   then  i2Rgb.red <= 737;
      elsif (i1Rgb.red   >= 740 and   i1Rgb.red <= (749+gain))   then  i2Rgb.red <= 747;
      elsif (i1Rgb.red   >= 750 and   i1Rgb.red <= (759+gain))   then  i2Rgb.red <= 757;
      elsif (i1Rgb.red   >= 760 and   i1Rgb.red <= (769+gain))   then  i2Rgb.red <= 767;
      elsif (i1Rgb.red   >= 770 and   i1Rgb.red <= (779+gain))   then  i2Rgb.red <= 777;
      elsif (i1Rgb.red   >= 780 and   i1Rgb.red <= (789+gain))   then  i2Rgb.red <= 787;
      elsif (i1Rgb.red   >= 790 and   i1Rgb.red <= (799+gain))   then  i2Rgb.red <= 797;
      elsif (i1Rgb.red   >= 800 and   i1Rgb.red <= (809+gain))   then  i2Rgb.red <= 807;
      elsif (i1Rgb.red   >= 810 and   i1Rgb.red <= (819+gain))   then  i2Rgb.red <= 817;
      elsif (i1Rgb.red   >= 820 and   i1Rgb.red <= (829+gain))   then  i2Rgb.red <= 827;
      elsif (i1Rgb.red   >= 830 and   i1Rgb.red <= (839+gain))   then  i2Rgb.red <= 837;
      elsif (i1Rgb.red   >= 840 and   i1Rgb.red <= (849+gain))   then  i2Rgb.red <= 847;
      elsif (i1Rgb.red   >= 850 and   i1Rgb.red <= (859+gain))   then  i2Rgb.red <= 857;
      elsif (i1Rgb.red   >= 860 and   i1Rgb.red <= (869+gain))   then  i2Rgb.red <= 867;
      elsif (i1Rgb.red   >= 870 and   i1Rgb.red <= (879+gain))   then  i2Rgb.red <= 877;
      elsif (i1Rgb.red   >= 880 and   i1Rgb.red <= (889+gain))   then  i2Rgb.red <= 887;
      elsif (i1Rgb.red   >= 890 and   i1Rgb.red <= (899+gain))   then  i2Rgb.red <= 897;
      elsif (i1Rgb.red   >= 900 and   i1Rgb.red <= (909+gain))   then  i2Rgb.red <= 907;
      elsif (i1Rgb.red   >= 910 and   i1Rgb.red <= (919+gain))   then  i2Rgb.red <= 917;
      elsif (i1Rgb.red   >= 920 and   i1Rgb.red <= (929+gain))   then  i2Rgb.red <= 927;
      elsif (i1Rgb.red   >= 930 and   i1Rgb.red <= (939+gain))   then  i2Rgb.red <= 937;
      elsif (i1Rgb.red   >= 940 and   i1Rgb.red <= (949+gain))   then  i2Rgb.red <= 947;
      elsif (i1Rgb.red   >= 950 and   i1Rgb.red <= (959+gain))   then  i2Rgb.red <= 957;
      elsif (i1Rgb.red   >= 960 and   i1Rgb.red <= (969+gain))   then  i2Rgb.red <= 967;
      elsif (i1Rgb.red   >= 970 and   i1Rgb.red <= (979+gain))   then  i2Rgb.red <= 977;
      elsif (i1Rgb.red   >= 980 and   i1Rgb.red <= (989+gain))   then  i2Rgb.red <= 987;
      elsif (i1Rgb.red   >= 990 and   i1Rgb.red <= (999+gain))   then  i2Rgb.red <= 997;
      elsif (i1Rgb.red   >= 1000 and  i1Rgb.red <= (1009+gain))  then  i2Rgb.red <= 1007;
      elsif (i1Rgb.red   >= 1010 and  i1Rgb.red <= (1019+gain))  then  i2Rgb.red <= 1017;
      elsif (i1Rgb.red   >= 1020 and  i1Rgb.red <= 1023)         then  i2Rgb.red <= 1023;
      else                                                       
        i2Rgb.red <= i1Rgb.red;
      end if;
    end if;
end process;
process (clk) begin
    if rising_edge(clk) then
      if (i1Rgb.green   >= 0 and     i1Rgb.green <= 9)               then  i2Rgb.green <= 7;
      elsif (i1Rgb.green   >= 10 and    i1Rgb.green <= (19))         then  i2Rgb.green <= 17;
      elsif (i1Rgb.green   >= 20 and    i1Rgb.green <= (29))         then  i2Rgb.green <= 27;
      elsif (i1Rgb.green   >= 30 and    i1Rgb.green <= (39+gain))    then  i2Rgb.green <= 37;
      elsif (i1Rgb.green   >= 40 and    i1Rgb.green <= (49+gain))    then  i2Rgb.green <= 47;
      elsif (i1Rgb.green   >= 50 and    i1Rgb.green <= (59+gain))    then  i2Rgb.green <= 57;
      elsif (i1Rgb.green   >= 60 and    i1Rgb.green <= (69+gain))    then  i2Rgb.green <= 67;
      elsif (i1Rgb.green   >= 70 and    i1Rgb.green <= (79+gain))    then  i2Rgb.green <= 77;
      elsif (i1Rgb.green   >= 80 and    i1Rgb.green <= (89+gain))    then  i2Rgb.green <= 87;
      elsif (i1Rgb.green   >= 90 and    i1Rgb.green <= (99+gain))    then  i2Rgb.green <= 97;
      elsif (i1Rgb.green   >= 100 and   i1Rgb.green <= (109+gain))   then  i2Rgb.green <= 107;
      elsif (i1Rgb.green   >= 110 and   i1Rgb.green <= (119+gain))   then  i2Rgb.green <= 117;
      elsif (i1Rgb.green   >= 120 and   i1Rgb.green <= (129+gain))   then  i2Rgb.green <= 127;
      elsif (i1Rgb.green   >= 130 and   i1Rgb.green <= (139+gain))   then  i2Rgb.green <= 137;
      elsif (i1Rgb.green   >= 140 and   i1Rgb.green <= (149+gain))   then  i2Rgb.green <= 147;
      elsif (i1Rgb.green   >= 150 and   i1Rgb.green <= (159+gain))   then  i2Rgb.green <= 157;
      elsif (i1Rgb.green   >= 160 and   i1Rgb.green <= (169+gain))   then  i2Rgb.green <= 167;
      elsif (i1Rgb.green   >= 170 and   i1Rgb.green <= (179+gain))   then  i2Rgb.green <= 177;
      elsif (i1Rgb.green   >= 180 and   i1Rgb.green <= (189+gain))   then  i2Rgb.green <= 187;
      elsif (i1Rgb.green   >= 190 and   i1Rgb.green <= (199+gain))   then  i2Rgb.green <= 197;
      elsif (i1Rgb.green   >= 200 and   i1Rgb.green <= (209+gain))   then  i2Rgb.green <= 207;
      elsif (i1Rgb.green   >= 210 and   i1Rgb.green <= (219+gain))   then  i2Rgb.green <= 217;
      elsif (i1Rgb.green   >= 220 and   i1Rgb.green <= (229+gain))   then  i2Rgb.green <= 227;
      elsif (i1Rgb.green   >= 230 and   i1Rgb.green <= (239+gain))   then  i2Rgb.green <= 237;
      elsif (i1Rgb.green   >= 240 and   i1Rgb.green <= (249+gain))   then  i2Rgb.green <= 247;
      elsif (i1Rgb.green   >= 250 and   i1Rgb.green <= (259+gain))   then  i2Rgb.green <= 257;
      elsif (i1Rgb.green   >= 260 and   i1Rgb.green <= (269+gain))   then  i2Rgb.green <= 267;
      elsif (i1Rgb.green   >= 270 and   i1Rgb.green <= (279+gain))   then  i2Rgb.green <= 277;
      elsif (i1Rgb.green   >= 280 and   i1Rgb.green <= (289+gain))   then  i2Rgb.green <= 287;
      elsif (i1Rgb.green   >= 290 and   i1Rgb.green <= (299+gain))   then  i2Rgb.green <= 297;
      elsif (i1Rgb.green   >= 300 and   i1Rgb.green <= (309+gain))   then  i2Rgb.green <= 307;
      elsif (i1Rgb.green   >= 310 and   i1Rgb.green <= (319+gain))   then  i2Rgb.green <= 317;
      elsif (i1Rgb.green   >= 320 and   i1Rgb.green <= (329+gain))   then  i2Rgb.green <= 327;
      elsif (i1Rgb.green   >= 330 and   i1Rgb.green <= (339+gain))   then  i2Rgb.green <= 337;
      elsif (i1Rgb.green   >= 340 and   i1Rgb.green <= (349+gain))   then  i2Rgb.green <= 347;
      elsif (i1Rgb.green   >= 350 and   i1Rgb.green <= (359+gain))   then  i2Rgb.green <= 357;
      elsif (i1Rgb.green   >= 360 and   i1Rgb.green <= (369+gain))   then  i2Rgb.green <= 367;
      elsif (i1Rgb.green   >= 370 and   i1Rgb.green <= (379+gain))   then  i2Rgb.green <= 377;
      elsif (i1Rgb.green   >= 380 and   i1Rgb.green <= (389+gain))   then  i2Rgb.green <= 387;
      elsif (i1Rgb.green   >= 390 and   i1Rgb.green <= (399+gain))   then  i2Rgb.green <= 397;
      elsif (i1Rgb.green   >= 400 and   i1Rgb.green <= (409+gain))   then  i2Rgb.green <= 407;
      elsif (i1Rgb.green   >= 400 and   i1Rgb.green <= (409+gain))   then  i2Rgb.green <= 407;
      elsif (i1Rgb.green   >= 410 and   i1Rgb.green <= (419+gain))   then  i2Rgb.green <= 417;
      elsif (i1Rgb.green   >= 420 and   i1Rgb.green <= (429+gain))   then  i2Rgb.green <= 427;
      elsif (i1Rgb.green   >= 430 and   i1Rgb.green <= (439+gain))   then  i2Rgb.green <= 437;
      elsif (i1Rgb.green   >= 440 and   i1Rgb.green <= (449+gain))   then  i2Rgb.green <= 447;
      elsif (i1Rgb.green   >= 450 and   i1Rgb.green <= (459+gain))   then  i2Rgb.green <= 457;
      elsif (i1Rgb.green   >= 460 and   i1Rgb.green <= (469+gain))   then  i2Rgb.green <= 467;
      elsif (i1Rgb.green   >= 470 and   i1Rgb.green <= (479+gain))   then  i2Rgb.green <= 477;
      elsif (i1Rgb.green   >= 480 and   i1Rgb.green <= (489+gain))   then  i2Rgb.green <= 487;
      elsif (i1Rgb.green   >= 490 and   i1Rgb.green <= (499+gain))   then  i2Rgb.green <= 497;
      elsif (i1Rgb.green   >= 500 and   i1Rgb.green <= (509+gain))   then  i2Rgb.green <= 507;
      elsif (i1Rgb.green   >= 510 and   i1Rgb.green <= (519+gain))   then  i2Rgb.green <= 517;
      elsif (i1Rgb.green   >= 520 and   i1Rgb.green <= (529+gain))   then  i2Rgb.green <= 527;
      elsif (i1Rgb.green   >= 530 and   i1Rgb.green <= (539+gain))   then  i2Rgb.green <= 537;
      elsif (i1Rgb.green   >= 540 and   i1Rgb.green <= (549+gain))   then  i2Rgb.green <= 547;
      elsif (i1Rgb.green   >= 550 and   i1Rgb.green <= (559+gain))   then  i2Rgb.green <= 557;
      elsif (i1Rgb.green   >= 560 and   i1Rgb.green <= (569+gain))   then  i2Rgb.green <= 567;
      elsif (i1Rgb.green   >= 570 and   i1Rgb.green <= (579+gain))   then  i2Rgb.green <= 577;
      elsif (i1Rgb.green   >= 580 and   i1Rgb.green <= (589+gain))   then  i2Rgb.green <= 587;
      elsif (i1Rgb.green   >= 590 and   i1Rgb.green <= (599+gain))   then  i2Rgb.green <= 597;
      elsif (i1Rgb.green   >= 600 and   i1Rgb.green <= (609+gain))   then  i2Rgb.green <= 607;
      elsif (i1Rgb.green   >= 610 and   i1Rgb.green <= (619+gain))   then  i2Rgb.green <= 617;
      elsif (i1Rgb.green   >= 620 and   i1Rgb.green <= (629+gain))   then  i2Rgb.green <= 627;
      elsif (i1Rgb.green   >= 630 and   i1Rgb.green <= (639+gain))   then  i2Rgb.green <= 637;
      elsif (i1Rgb.green   >= 640 and   i1Rgb.green <= (649+gain))   then  i2Rgb.green <= 647;
      elsif (i1Rgb.green   >= 650 and   i1Rgb.green <= (659+gain))   then  i2Rgb.green <= 657;
      elsif (i1Rgb.green   >= 660 and   i1Rgb.green <= (669+gain))   then  i2Rgb.green <= 667;
      elsif (i1Rgb.green   >= 670 and   i1Rgb.green <= (679+gain))   then  i2Rgb.green <= 677;
      elsif (i1Rgb.green   >= 680 and   i1Rgb.green <= (689+gain))   then  i2Rgb.green <= 687;
      elsif (i1Rgb.green   >= 690 and   i1Rgb.green <= (699+gain))   then  i2Rgb.green <= 697;
      elsif (i1Rgb.green   >= 700 and   i1Rgb.green <= (709+gain))   then  i2Rgb.green <= 707;
      elsif (i1Rgb.green   >= 710 and   i1Rgb.green <= (719+gain))   then  i2Rgb.green <= 717;
      elsif (i1Rgb.green   >= 720 and   i1Rgb.green <= (729+gain))   then  i2Rgb.green <= 727;
      elsif (i1Rgb.green   >= 730 and   i1Rgb.green <= (739+gain))   then  i2Rgb.green <= 737;
      elsif (i1Rgb.green   >= 740 and   i1Rgb.green <= (749+gain))   then  i2Rgb.green <= 747;
      elsif (i1Rgb.green   >= 750 and   i1Rgb.green <= (759+gain))   then  i2Rgb.green <= 757;
      elsif (i1Rgb.green   >= 760 and   i1Rgb.green <= (769+gain))   then  i2Rgb.green <= 767;
      elsif (i1Rgb.green   >= 770 and   i1Rgb.green <= (779+gain))   then  i2Rgb.green <= 777;
      elsif (i1Rgb.green   >= 780 and   i1Rgb.green <= (789+gain))   then  i2Rgb.green <= 787;
      elsif (i1Rgb.green   >= 790 and   i1Rgb.green <= (799+gain))   then  i2Rgb.green <= 797;
      elsif (i1Rgb.green   >= 800 and   i1Rgb.green <= (809+gain))   then  i2Rgb.green <= 807;
      elsif (i1Rgb.green   >= 810 and   i1Rgb.green <= (819+gain))   then  i2Rgb.green <= 817;
      elsif (i1Rgb.green   >= 820 and   i1Rgb.green <= (829+gain))   then  i2Rgb.green <= 827;
      elsif (i1Rgb.green   >= 830 and   i1Rgb.green <= (839+gain))   then  i2Rgb.green <= 837;
      elsif (i1Rgb.green   >= 840 and   i1Rgb.green <= (849+gain))   then  i2Rgb.green <= 847;
      elsif (i1Rgb.green   >= 850 and   i1Rgb.green <= (859+gain))   then  i2Rgb.green <= 857;
      elsif (i1Rgb.green   >= 860 and   i1Rgb.green <= (869+gain))   then  i2Rgb.green <= 867;
      elsif (i1Rgb.green   >= 870 and   i1Rgb.green <= (879+gain))   then  i2Rgb.green <= 877;
      elsif (i1Rgb.green   >= 880 and   i1Rgb.green <= (889+gain))   then  i2Rgb.green <= 887;
      elsif (i1Rgb.green   >= 890 and   i1Rgb.green <= (899+gain))   then  i2Rgb.green <= 897;
      elsif (i1Rgb.green   >= 900 and   i1Rgb.green <= (909+gain))   then  i2Rgb.green <= 907;
      elsif (i1Rgb.green   >= 910 and   i1Rgb.green <= (919+gain))   then  i2Rgb.green <= 917;
      elsif (i1Rgb.green   >= 920 and   i1Rgb.green <= (929+gain))   then  i2Rgb.green <= 927;
      elsif (i1Rgb.green   >= 930 and   i1Rgb.green <= (939+gain))   then  i2Rgb.green <= 937;
      elsif (i1Rgb.green   >= 940 and   i1Rgb.green <= (949+gain))   then  i2Rgb.green <= 947;
      elsif (i1Rgb.green   >= 950 and   i1Rgb.green <= (959+gain))   then  i2Rgb.green <= 957;
      elsif (i1Rgb.green   >= 960 and   i1Rgb.green <= (969+gain))   then  i2Rgb.green <= 967;
      elsif (i1Rgb.green   >= 970 and   i1Rgb.green <= (979+gain))   then  i2Rgb.green <= 977;
      elsif (i1Rgb.green   >= 980 and   i1Rgb.green <= (989+gain))   then  i2Rgb.green <= 987;
      elsif (i1Rgb.green   >= 990 and   i1Rgb.green <= (999+gain))   then  i2Rgb.green <= 997;
      elsif (i1Rgb.green   >= 1000 and  i1Rgb.green <= (1009+gain))  then  i2Rgb.green <= 1007;
      elsif (i1Rgb.green   >= 1010 and  i1Rgb.green <= (1019+gain))  then  i2Rgb.green <= 1017;
      elsif (i1Rgb.green   >= 1020 and  i1Rgb.green <= 1023)         then  i2Rgb.green <= 1023;
      else                                                       
        i2Rgb.green <= i1Rgb.green;
      end if;
    end if;
end process;
process (clk) begin
    if rising_edge(clk) then
      if (i1Rgb.blue   >= 0 and     i1Rgb.blue <= 9)               then  i2Rgb.blue <= 7;
      elsif (i1Rgb.blue   >= 10 and    i1Rgb.blue <= (19))         then  i2Rgb.blue <= 17;
      elsif (i1Rgb.blue   >= 20 and    i1Rgb.blue <= (29))         then  i2Rgb.blue <= 27;
      elsif (i1Rgb.blue   >= 30 and    i1Rgb.blue <= (39+gain))    then  i2Rgb.blue <= 37;
      elsif (i1Rgb.blue   >= 40 and    i1Rgb.blue <= (49+gain))    then  i2Rgb.blue <= 47;
      elsif (i1Rgb.blue   >= 50 and    i1Rgb.blue <= (59+gain))    then  i2Rgb.blue <= 57;
      elsif (i1Rgb.blue   >= 60 and    i1Rgb.blue <= (69+gain))    then  i2Rgb.blue <= 67;
      elsif (i1Rgb.blue   >= 70 and    i1Rgb.blue <= (79+gain))    then  i2Rgb.blue <= 77;
      elsif (i1Rgb.blue   >= 80 and    i1Rgb.blue <= (89+gain))    then  i2Rgb.blue <= 87;
      elsif (i1Rgb.blue   >= 90 and    i1Rgb.blue <= (99+gain))    then  i2Rgb.blue <= 97;
      elsif (i1Rgb.blue   >= 100 and   i1Rgb.blue <= (109+gain))   then  i2Rgb.blue <= 107;
      elsif (i1Rgb.blue   >= 110 and   i1Rgb.blue <= (119+gain))   then  i2Rgb.blue <= 117;
      elsif (i1Rgb.blue   >= 120 and   i1Rgb.blue <= (129+gain))   then  i2Rgb.blue <= 127;
      elsif (i1Rgb.blue   >= 130 and   i1Rgb.blue <= (139+gain))   then  i2Rgb.blue <= 137;
      elsif (i1Rgb.blue   >= 140 and   i1Rgb.blue <= (149+gain))   then  i2Rgb.blue <= 147;
      elsif (i1Rgb.blue   >= 150 and   i1Rgb.blue <= (159+gain))   then  i2Rgb.blue <= 157;
      elsif (i1Rgb.blue   >= 160 and   i1Rgb.blue <= (169+gain))   then  i2Rgb.blue <= 167;
      elsif (i1Rgb.blue   >= 170 and   i1Rgb.blue <= (179+gain))   then  i2Rgb.blue <= 177;
      elsif (i1Rgb.blue   >= 180 and   i1Rgb.blue <= (189+gain))   then  i2Rgb.blue <= 187;
      elsif (i1Rgb.blue   >= 190 and   i1Rgb.blue <= (199+gain))   then  i2Rgb.blue <= 197;
      elsif (i1Rgb.blue   >= 200 and   i1Rgb.blue <= (209+gain))   then  i2Rgb.blue <= 207;
      elsif (i1Rgb.blue   >= 210 and   i1Rgb.blue <= (219+gain))   then  i2Rgb.blue <= 217;
      elsif (i1Rgb.blue   >= 220 and   i1Rgb.blue <= (229+gain))   then  i2Rgb.blue <= 227;
      elsif (i1Rgb.blue   >= 230 and   i1Rgb.blue <= (239+gain))   then  i2Rgb.blue <= 237;
      elsif (i1Rgb.blue   >= 240 and   i1Rgb.blue <= (249+gain))   then  i2Rgb.blue <= 247;
      elsif (i1Rgb.blue   >= 250 and   i1Rgb.blue <= (259+gain))   then  i2Rgb.blue <= 257;
      elsif (i1Rgb.blue   >= 260 and   i1Rgb.blue <= (269+gain))   then  i2Rgb.blue <= 267;
      elsif (i1Rgb.blue   >= 270 and   i1Rgb.blue <= (279+gain))   then  i2Rgb.blue <= 277;
      elsif (i1Rgb.blue   >= 280 and   i1Rgb.blue <= (289+gain))   then  i2Rgb.blue <= 287;
      elsif (i1Rgb.blue   >= 290 and   i1Rgb.blue <= (299+gain))   then  i2Rgb.blue <= 297;
      elsif (i1Rgb.blue   >= 300 and   i1Rgb.blue <= (309+gain))   then  i2Rgb.blue <= 307;
      elsif (i1Rgb.blue   >= 310 and   i1Rgb.blue <= (319+gain))   then  i2Rgb.blue <= 317;
      elsif (i1Rgb.blue   >= 320 and   i1Rgb.blue <= (329+gain))   then  i2Rgb.blue <= 327;
      elsif (i1Rgb.blue   >= 330 and   i1Rgb.blue <= (339+gain))   then  i2Rgb.blue <= 337;
      elsif (i1Rgb.blue   >= 340 and   i1Rgb.blue <= (349+gain))   then  i2Rgb.blue <= 347;
      elsif (i1Rgb.blue   >= 350 and   i1Rgb.blue <= (359+gain))   then  i2Rgb.blue <= 357;
      elsif (i1Rgb.blue   >= 360 and   i1Rgb.blue <= (369+gain))   then  i2Rgb.blue <= 367;
      elsif (i1Rgb.blue   >= 370 and   i1Rgb.blue <= (379+gain))   then  i2Rgb.blue <= 377;
      elsif (i1Rgb.blue   >= 380 and   i1Rgb.blue <= (389+gain))   then  i2Rgb.blue <= 387;
      elsif (i1Rgb.blue   >= 390 and   i1Rgb.blue <= (399+gain))   then  i2Rgb.blue <= 397;
      elsif (i1Rgb.blue   >= 400 and   i1Rgb.blue <= (409+gain))   then  i2Rgb.blue <= 407;
      elsif (i1Rgb.blue   >= 400 and   i1Rgb.blue <= (409+gain))   then  i2Rgb.blue <= 407;
      elsif (i1Rgb.blue   >= 410 and   i1Rgb.blue <= (419+gain))   then  i2Rgb.blue <= 417;
      elsif (i1Rgb.blue   >= 420 and   i1Rgb.blue <= (429+gain))   then  i2Rgb.blue <= 427;
      elsif (i1Rgb.blue   >= 430 and   i1Rgb.blue <= (439+gain))   then  i2Rgb.blue <= 437;
      elsif (i1Rgb.blue   >= 440 and   i1Rgb.blue <= (449+gain))   then  i2Rgb.blue <= 447;
      elsif (i1Rgb.blue   >= 450 and   i1Rgb.blue <= (459+gain))   then  i2Rgb.blue <= 457;
      elsif (i1Rgb.blue   >= 460 and   i1Rgb.blue <= (469+gain))   then  i2Rgb.blue <= 467;
      elsif (i1Rgb.blue   >= 470 and   i1Rgb.blue <= (479+gain))   then  i2Rgb.blue <= 477;
      elsif (i1Rgb.blue   >= 480 and   i1Rgb.blue <= (489+gain))   then  i2Rgb.blue <= 487;
      elsif (i1Rgb.blue   >= 490 and   i1Rgb.blue <= (499+gain))   then  i2Rgb.blue <= 497;
      elsif (i1Rgb.blue   >= 500 and   i1Rgb.blue <= (509+gain))   then  i2Rgb.blue <= 507;
      elsif (i1Rgb.blue   >= 510 and   i1Rgb.blue <= (519+gain))   then  i2Rgb.blue <= 517;
      elsif (i1Rgb.blue   >= 520 and   i1Rgb.blue <= (529+gain))   then  i2Rgb.blue <= 527;
      elsif (i1Rgb.blue   >= 530 and   i1Rgb.blue <= (539+gain))   then  i2Rgb.blue <= 537;
      elsif (i1Rgb.blue   >= 540 and   i1Rgb.blue <= (549+gain))   then  i2Rgb.blue <= 547;
      elsif (i1Rgb.blue   >= 550 and   i1Rgb.blue <= (559+gain))   then  i2Rgb.blue <= 557;
      elsif (i1Rgb.blue   >= 560 and   i1Rgb.blue <= (569+gain))   then  i2Rgb.blue <= 567;
      elsif (i1Rgb.blue   >= 570 and   i1Rgb.blue <= (579+gain))   then  i2Rgb.blue <= 577;
      elsif (i1Rgb.blue   >= 580 and   i1Rgb.blue <= (589+gain))   then  i2Rgb.blue <= 587;
      elsif (i1Rgb.blue   >= 590 and   i1Rgb.blue <= (599+gain))   then  i2Rgb.blue <= 597;
      elsif (i1Rgb.blue   >= 600 and   i1Rgb.blue <= (609+gain))   then  i2Rgb.blue <= 607;
      elsif (i1Rgb.blue   >= 610 and   i1Rgb.blue <= (619+gain))   then  i2Rgb.blue <= 617;
      elsif (i1Rgb.blue   >= 620 and   i1Rgb.blue <= (629+gain))   then  i2Rgb.blue <= 627;
      elsif (i1Rgb.blue   >= 630 and   i1Rgb.blue <= (639+gain))   then  i2Rgb.blue <= 637;
      elsif (i1Rgb.blue   >= 640 and   i1Rgb.blue <= (649+gain))   then  i2Rgb.blue <= 647;
      elsif (i1Rgb.blue   >= 650 and   i1Rgb.blue <= (659+gain))   then  i2Rgb.blue <= 657;
      elsif (i1Rgb.blue   >= 660 and   i1Rgb.blue <= (669+gain))   then  i2Rgb.blue <= 667;
      elsif (i1Rgb.blue   >= 670 and   i1Rgb.blue <= (679+gain))   then  i2Rgb.blue <= 677;
      elsif (i1Rgb.blue   >= 680 and   i1Rgb.blue <= (689+gain))   then  i2Rgb.blue <= 687;
      elsif (i1Rgb.blue   >= 690 and   i1Rgb.blue <= (699+gain))   then  i2Rgb.blue <= 697;
      elsif (i1Rgb.blue   >= 700 and   i1Rgb.blue <= (709+gain))   then  i2Rgb.blue <= 707;
      elsif (i1Rgb.blue   >= 710 and   i1Rgb.blue <= (719+gain))   then  i2Rgb.blue <= 717;
      elsif (i1Rgb.blue   >= 720 and   i1Rgb.blue <= (729+gain))   then  i2Rgb.blue <= 727;
      elsif (i1Rgb.blue   >= 730 and   i1Rgb.blue <= (739+gain))   then  i2Rgb.blue <= 737;
      elsif (i1Rgb.blue   >= 740 and   i1Rgb.blue <= (749+gain))   then  i2Rgb.blue <= 747;
      elsif (i1Rgb.blue   >= 750 and   i1Rgb.blue <= (759+gain))   then  i2Rgb.blue <= 757;
      elsif (i1Rgb.blue   >= 760 and   i1Rgb.blue <= (769+gain))   then  i2Rgb.blue <= 767;
      elsif (i1Rgb.blue   >= 770 and   i1Rgb.blue <= (779+gain))   then  i2Rgb.blue <= 777;
      elsif (i1Rgb.blue   >= 780 and   i1Rgb.blue <= (789+gain))   then  i2Rgb.blue <= 787;
      elsif (i1Rgb.blue   >= 790 and   i1Rgb.blue <= (799+gain))   then  i2Rgb.blue <= 797;
      elsif (i1Rgb.blue   >= 800 and   i1Rgb.blue <= (809+gain))   then  i2Rgb.blue <= 807;
      elsif (i1Rgb.blue   >= 810 and   i1Rgb.blue <= (819+gain))   then  i2Rgb.blue <= 817;
      elsif (i1Rgb.blue   >= 820 and   i1Rgb.blue <= (829+gain))   then  i2Rgb.blue <= 827;
      elsif (i1Rgb.blue   >= 830 and   i1Rgb.blue <= (839+gain))   then  i2Rgb.blue <= 837;
      elsif (i1Rgb.blue   >= 840 and   i1Rgb.blue <= (849+gain))   then  i2Rgb.blue <= 847;
      elsif (i1Rgb.blue   >= 850 and   i1Rgb.blue <= (859+gain))   then  i2Rgb.blue <= 857;
      elsif (i1Rgb.blue   >= 860 and   i1Rgb.blue <= (869+gain))   then  i2Rgb.blue <= 867;
      elsif (i1Rgb.blue   >= 870 and   i1Rgb.blue <= (879+gain))   then  i2Rgb.blue <= 877;
      elsif (i1Rgb.blue   >= 880 and   i1Rgb.blue <= (889+gain))   then  i2Rgb.blue <= 887;
      elsif (i1Rgb.blue   >= 890 and   i1Rgb.blue <= (899+gain))   then  i2Rgb.blue <= 897;
      elsif (i1Rgb.blue   >= 900 and   i1Rgb.blue <= (909+gain))   then  i2Rgb.blue <= 907;
      elsif (i1Rgb.blue   >= 910 and   i1Rgb.blue <= (919+gain))   then  i2Rgb.blue <= 917;
      elsif (i1Rgb.blue   >= 920 and   i1Rgb.blue <= (929+gain))   then  i2Rgb.blue <= 927;
      elsif (i1Rgb.blue   >= 930 and   i1Rgb.blue <= (939+gain))   then  i2Rgb.blue <= 937;
      elsif (i1Rgb.blue   >= 940 and   i1Rgb.blue <= (949+gain))   then  i2Rgb.blue <= 947;
      elsif (i1Rgb.blue   >= 950 and   i1Rgb.blue <= (959+gain))   then  i2Rgb.blue <= 957;
      elsif (i1Rgb.blue   >= 960 and   i1Rgb.blue <= (969+gain))   then  i2Rgb.blue <= 967;
      elsif (i1Rgb.blue   >= 970 and   i1Rgb.blue <= (979+gain))   then  i2Rgb.blue <= 977;
      elsif (i1Rgb.blue   >= 980 and   i1Rgb.blue <= (989+gain))   then  i2Rgb.blue <= 987;
      elsif (i1Rgb.blue   >= 990 and   i1Rgb.blue <= (999+gain))   then  i2Rgb.blue <= 997;
      elsif (i1Rgb.blue   >= 1000 and  i1Rgb.blue <= (1009+gain))  then  i2Rgb.blue <= 1007;
      elsif (i1Rgb.blue   >= 1010 and  i1Rgb.blue <= (1019+gain))  then  i2Rgb.blue <= 1017;
      elsif (i1Rgb.blue   >= 1020 and  i1Rgb.blue <= 1023)         then  i2Rgb.blue <= 1023;
      else                                                       
        i2Rgb.blue <= i1Rgb.blue;
      end if;
    end if;
end process;
 oRgb.red   <= std_logic_vector(to_unsigned(i2Rgb.red, 10));
 oRgb.green <= std_logic_vector(to_unsigned(i2Rgb.green, 10));
 oRgb.blue  <= std_logic_vector(to_unsigned(i2Rgb.blue, 10));
 oRgb.valid <= i1Rgb.valid;
 oRgb.eol   <= rgbSyncEol;
 oRgb.sof   <= rgbSyncSof;
 oRgb.eof   <= rgbSyncEof;
end Behavioral;